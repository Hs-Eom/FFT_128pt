library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Mult is
    generic(BW : integer := 16;
            N : integer := 64
    );
    port(
        cnt : in std_logic_vector(5 downto 0);
        In_Real, In_Imag : in std_logic_vector(BW downto 0);

        Out_Real, Out_Imag : out std_logic_vector(BW downto 0)
    );
end Mult;

architecture rtl of Mult is
    --12bit in array of 64
    subtype bit12 is std_logic_vector(11 downto 0);
    type bit12_arr64 is array(0 to 63) of bit12;

    signal W_tmp_re, W_tmp_im : bit12;

    signal buf_re0, buf_im0 : signed(BW +13 downto 0);
    signal buf_re1, buf_im1 : signed(BW +13 downto 0);
    signal buf_re  : signed(BW +13 downto 0);
    signal buf_im  : signed(BW+13 downto 0);   
    signal cnt_num : integer;

    --Twiddle Factors
    constant W_re : bit12_arr64 :=(
    "010000000000", "001111111110", "001111111011", "001111110100",
    "001111101100", "001111100001", "001111010011", "001111000100",
    "001110110010", "001110011101", "001110000111", "001101101110",
    "001101010011", "001100110110", "001100010111", "001011110110",
    "001011010100", "001010101111", "001010001001", "001001100001",
    "001000111000", "001000001110", "000111100010", "000110110101",
    "000110000111", "000101011000", "000100101001", "000011111000",
    "000011000111", "000010010110", "000001100100", "000000110010",
    "000000000000", "111111001101", "111110011011", "111101101001",
    "111100111000", "111100000111", "111011010110", "111010100111",
    "111001111000", "111001001010", "111000011101", "110111110001",
    "110111000111", "110110011110", "110101110110", "110101010000",
    "110100101011", "110100001001", "110011101000", "110011001001",
    "110010101100", "110010010001", "110001111000", "110001100010",
    "110001001101", "110000111011", "110000101100", "110000011110",
    "110000010011", "110000001011", "110000000100", "110000000001"
    );
    constant W_im : bit12_arr64 := (
    "000000000000", "111111001101", "111110011011", "111101101001",
    "111100111000", "111100000111", "111011010110", "111010100111",
    "111001111000", "111001001010", "111000011101", "110111110001",
    "110111000111", "110110011110", "110101110110", "110101010000",
    "110100101011", "110100001001", "110011101000", "110011001001",
    "110010101100", "110010010001", "110001111000", "110001100010",
    "110001001101", "110000111011", "110000101100", "110000011110",
    "110000010011", "110000001011", "110000000100", "110000000001",
    "110000000000", "110000000001", "110000000100", "110000001011",
    "110000010011", "110000011110", "110000101100", "110000111011",
    "110001001101", "110001100010", "110001111000", "110010010001",
    "110010101100", "110011001001", "110011101000", "110100001001",
    "110100101011", "110101010000", "110101110110", "110110011110",
    "110111000111", "110111110001", "111000011101", "111001001010",
    "111001111000", "111010100111", "111011010110", "111100000111",
    "111100111000", "111101101001", "111110011011", "111111001101"
    );

    begin
        W_tmp_re <= W_re(to_integer(unsigned(cnt)));
        W_tmp_im <= W_im(to_integer(unsigned(cnt)));

        buf_re0 <= resize(signed(In_Real) * signed(W_tmp_re),BW+14); --(29:0) BW+13 = (BW+1)+12
        buf_re1 <= resize(signed(In_Imag) * signed(W_tmp_im),BW+14);
        buf_im0 <= resize(signed(In_Real) * signed(W_tmp_im),BW+14);
        buf_im1 <= resize(signed(In_Imag) * signed(W_tmp_re),BW+14);

        buf_re <= signed(buf_re0 - buf_re1);
        buf_im <= signed(buf_im0 + buf_im1);


        Out_Real <= std_logic_vector(buf_re(BW + 13) & buf_re(BW + 9 downto 10));
        Out_Imag <= std_logic_vector(buf_im(BW + 13) & buf_im(BW + 9 downto 10));

    end rtl;

